`timescale 1ns / 1ps

module qmult #(
	parameter Q = 15,
	parameter N = 32
)(
	 input	[N-1:0]	    i_multiplicand,
	 input	[N-1:0]   	i_multiplier  ,
	 output	[2*N-1:0]	r_result
	 //output	reg				ovr
);

assign r_result = $signed(i_multiplicand) * $signed(i_multiplier) ;
	 
//	The underlying assumption, here, is that both fixed-point values are of the same length (N,Q)
//		Because of this, the results will be of length N+N = 2N bits....
//		This also simplifies the hand-back of results, as the binimal point 
//		will always be in the same location...
	
//reg [2*N-1:0]	r_result;	//	Multiplication by 2 values of N bits requires a 
                            //		register that is N+N = 2N deep...
//reg [N-1:0]		r_RetVal;
	
//--------------------------------------------------------------------------------
//	assign o_result = r_RetVal;	//	Only handing back the same number of bits as we received...
											//		with fixed point in same location...
	
//---------------------------------------------------------------------------------
// always @(*)	begin						//	Do the multiply any time the inputs change
// 	r_result <= i_multiplicand[N-2:0] * i_multiplier[N-2:0];	//	removing the sign bits from the multiply - that 
// end															//	would introduce *big* errors	
//	ovr <= 1'b0;												//	reset overflow flag to zero
		
	
//	This always block will throw a warning, as it uses a & b, but only acts on changes in result...
//	always @(r_result) begin										// any time the result changes, we need to recompute the sign bit,
//		r_RetVal[N-1] <= i_multiplicand[N-1] ^ i_multiplier[N-1];	//		which is the XOR of the input sign bits...  (you do the truth table...)
//		r_RetVal[N-2:0] <= r_result[N-2+Q:Q];						// and we also need to push the proper N bits of result up to 
//																	//		the calling entity...
//		if (r_result[2*N-2:N-1+Q] > 0)								// and finally, we need to check for an overflow
//			ovr <= 1'b1;
//		end

endmodule
